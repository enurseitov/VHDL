`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:36:08 09/12/2016 
// Design Name: 
// Module Name:    fourBitAdder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fourBitAdder(
    input [0:3] inA,
    input [0:3] inB,
    output [0:3] Result,
    output CarryOut,
    input CarryIn
    );


endmodule
